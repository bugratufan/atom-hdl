
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity $entity_name is
    port (
        i_clk : std_logic;
        i_rst : std_logic
    );
end entity;



architecture arch of $entity_name is
begin

end architecture;
