-- ===============================================================================================
-- (C) COPYRIGHT $year Rohde & Schwarz
-- All rights reserved.
-- ===============================================================================================
-- Creator: $pc_name
-- ===============================================================================================
-- Project           : $entity_name
-- File ID           : $file_name
-- Design Unit Name  :
-- Description       :
-- Comments          :
-- Revision          : %%
-- Last Changed Date : %%
-- Last Changed By   : %%
-- Designer
--          Name     : Bugra Tufan
--          E-mail   : btufan21@ku.edu.tr
-- ===============================================================================================
